timeunit 1s;

module test;
endmodule